-- emp_project_decl for the Phase-2 GT prototype
--
-- Defines constants for the whole project
--
library IEEE;
use IEEE.STD_LOGIC_1164.all;

use work.emp_framework_decl.all;
use work.emp_device_types.all;

-------------------------------------------------------------------------------
package emp_project_decl is

  constant PAYLOAD_REV : std_logic_vector(31 downto 0) := X"12345678";

  -- Latency buffer size
  constant LB_ADDR_WIDTH : integer := 10;

  -- Clock setup
  constant CLOCK_COMMON_RATIO : integer               := 36;
  constant CLOCK_RATIO        : integer               := 9;
  constant CLOCK_AUX_DIV      : clock_divisor_array_t := (36, 6, 3); -- 40 MHz, 240 MHz, 480 MHz

  constant ALGO_REPLICATION_IN_SRL : natural := 2;
  constant NUM_SLR                 : natural := 3;

  constant REGION_CONF : region_conf_array_t := (
    0  => (gty25, buf, no_fmt, buf, gty25),
    1  => (gty25, buf, no_fmt, buf, gty25),
    2  => (gty25, buf, no_fmt, buf, gty25),
    3  => (gty25, buf, no_fmt, buf, gty25),
    4  => kDummyRegion, -- HighSpeedBus
    5  => kDummyRegion, -- PCIe, AXI & TCDS
    6  => (gty25, buf, no_fmt, buf, gty25),
    7  => (gty25, buf, no_fmt, buf, gty25),
    8  => (gty25, buf, no_fmt, buf, gty25),
    9  => (gty25, buf, no_fmt, buf, gty25),
    10 => (gty25, buf, no_fmt, buf, gty25),
    11 => (gty25, buf, no_fmt, buf, gty25),
    12 => (gty25, buf, no_fmt, buf, gty25),
    13 => (gty25, buf, no_fmt, buf, gty25),
    14 => (gty25, buf, no_fmt, buf, gty25),
    -- Cross-chip
    15     => (gty25, buf, no_fmt, buf, gty25),
    16     => (gty25, buf, no_fmt, buf, gty25),
    17     => (gty25, buf, no_fmt, buf, gty25),
    18     => (gty25, buf, no_fmt, buf, gty25),
    19     => (gty25, buf, no_fmt, buf, gty25),
    20     => (gty25, buf, no_fmt, buf, gty25),
    21     => (gty25, buf, no_fmt, buf, gty25),
    22     => (gty25, buf, no_fmt, buf, gty25),
    23     => (gty25, buf, no_fmt, buf, gty25),
    24     => kDummyRegion, -- Unconnected
    25     => kDummyRegion, -- HighSpeedBus
    26     => (gty25, buf, no_fmt, buf, gty25),
    27     => (gty25, buf, no_fmt, buf, gty25),
    28     => (gty25, buf, no_fmt, buf, gty25),
    29     => (gty25, buf, no_fmt, buf, gty25),
    others => kDummyRegion
  );

end emp_project_decl;

-------------------------------------------------------------------------------

